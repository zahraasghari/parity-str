library ieee;
use ieee.std_logic_1164.all;

entity parity1 is

 port (a:in std_logic_vector(15 downto 0); 
     b:OUT std_logic
	);
	 end parity1 ;
	 
	 	 
	architecture logic of parity1 is
	
	begin
	b<=(a(0) xor a(1) xor a(2) xor a(3) xor a(4) xor a(5) xor a(6) xor a(7) xor a(8) xor a(9) xor a(10) xor a(11) xor a(12) xor a(13) xor a(14) xor a(15));
	
	 end architecture ;
